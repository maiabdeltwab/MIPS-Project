`timescale 1ns / 1ps

//
// 3rd year -Computer and Systems Engineering-
// Fayoum University
// Microprocessors (301)
// Pipelined Mips 32-bit project
// ____Group1____ 
// Supervised by: Dr.Mohammed Ibrahim
//


//pc reset to 00000000

module MIPS(
		input clk,
		input reset_b
    );
	 
	 
	 
	 //============================================ IF stage =============================================
	 wire [31:0] pc_new ,pc_new1 , pc_new2 , pc_new3 , pc_new4 , pc_new5 , pc_new6 ;
	 wire[31:0] pc_if;
	 reg pc_en_id;
	 
	Register 
	 #(
	 .WIDTH(32)
	 )
	 PC
	 (
	 .din(pc_new),
	 .dout(pc_if),
	 .en(pc_en_id),
	 .clk(clk),
	 .reset_b(reset_b)
	 );

	
	 wire[31:0] read_instr_if;
	 wire[31:0] instr_if;
	 reg if_id_enable;
	 
	 IMem IM(
	 .address(pc_if),
	 .dout(read_instr_if),
	 .enable(if_id_enable),
	 .clk(clk)
	 );
	 
	 
	 //if reset, the read instruction is nop
	 assign instr_if = (reset_b==0) ? 0 : read_instr_if;
	 
	 wire[31:0] pc_add_4_if;
	 wire[31:0] pc_add_1_if;
	 
	 assign pc_add_4_if= (reset_b==0) ? 0 : (pc_if+4);
	 assign pc_add_1_if= (reset_b==0) ? 0 : (pc_if+1);
	 
	 //PC select multiplexers
	 reg[31:0] pc_branch_mem , pc_jump_mem , pc_jumpr_mem ;


	wire  beq_sel_mem, bne_sel_mem, bgtz_sel_mem, blez_sel_mem, bgez_sel_mem, jump_sel_mem, jumpr_sel_mem ;
	
	assign pc_new1 =( beq_sel_mem==0 ) ? pc_add_4_if : pc_branch_mem;						// Branch IF Equal
	
	assign pc_new2 =( bne_sel_mem ==0 ) ?  pc_new1 : pc_branch_mem;							// Branch IF not Equal
	
	assign pc_new3 =( bgtz_sel_mem ==0 ) ?  pc_new2 : pc_branch_mem;							// Branch IF Bigger than (Bigger than zero)
	
	assign pc_new4 =( blez_sel_mem ==0 ) ?  pc_new3 : pc_branch_mem;							// Branch IF less than or Equal zero
	
	assign pc_new5 =( bgez_sel_mem ==0 ) ?  pc_new4 : pc_branch_mem;							// Branch IF Bigger than or Equal zero
	
	assign pc_new6 =( jump_sel_mem ==0 ) ?  pc_new5 : pc_jump_mem;							// Jump or Jump And Link
	
	assign pc_new =( jumpr_sel_mem ==0 ) ?  pc_new6 : pc_jumpr_mem;							// Jump Register | J A L R
	
	
	 
	 //====================================================ID stage============================================
	 
	 reg[31:0] pc_add_4_id;
	 reg[31:0] pc_add_1_id;
	 reg[31:0] instr_id;
	 
	 
	 
	 //IF/ID pipeline register
	 always @(posedge clk)
	 begin
		if(if_id_enable==1)
		begin
			pc_add_4_id <= pc_add_4_if;
			pc_add_1_id <= pc_add_1_if;
			instr_id <= instr_if;
		end
	end

	wire[4:0] rs_id,rt_id,rd_id,shamt_id;
	wire[5:0] opcode_id,func_id;
	wire[25:0] jumpConst_id;
	wire[15:0] imm16_id;
	
	assign rs_id=instr_id[25:21];
	assign rt_id=instr_id[20:16];
	assign rd_id=instr_id[15:11];
	assign shamt_id=instr_id[10:6];
	assign opcode_id=instr_id[31:26];
	assign func_id=instr_id[5:0];
	assign jumpConst_id=instr_id[25:0];
	assign imm16_id = instr_id[15:0];

	reg[4:0] rd_actual_wb;//register write index (from WB stage)
	wire[31:0] reg_wr_wb; //register 
	
	wire[31:0] reg_rd1_ex,reg_rd2_ex;
	
	
	reg id_ex_enable;
	
	reg regWrite_wb;//register file write control signal


	// hi and lo registers
	 reg lo_en_id;
	 reg hi_en_id;
	 
	 wire [31:0] lo_dataIn_wb;
	 wire [31:0] hi_dataIn_wb;	 
	 wire[31:0] lo_dataOut_id;
	 wire[31:0] hi_dataOut_id;	 

	 Register 
	 #(
	 .WIDTH(32)
	 )
	 lo
	 (
	 .din(lo_dataIn_wb),
	 .dout(lo_dataOut_id),
	 .en(lo_en_id),
	 .clk(clk),
	 .reset_b(reset_b)	 
	 );

	 Register 
	 #(
	 .WIDTH(32)
	 )
	 hi
	 (
	 .din(hi_dataIn_wb),
	 .dout(hi_dataOut_id),
	 .en(hi_en_id),
	 .clk(clk),
	 .reset_b(reset_b)	 
	 );


	
	RegFile RegFile(
		.rd1_index(rs_id),
		.rd2_index(rt_id),
		.wr_index(rd_actual_wb),
		.rd1_out(reg_rd1_ex),
		.rd2_out(reg_rd2_ex),
		.wr_in(reg_wr_wb),
		.regWrite(regWrite_wb),
		.regRead(id_ex_enable),
		.clk(clk)
	);
	
	wire regWrite_id;//generated by control but not used now    reg file write enable
	wire regDst_id; //selector for the write register source (0--> rt or 1--> rd) 
	wire aluSrc_id; //alu second operand source register 0--> from register file 1-->sign extended word
	wire beq_id;
	wire bne_id;
	wire blez_id;
	wire bgez_id;
	wire bgtz_id;
	wire jal_id;
	wire jr_id;
	wire j_id;
	wire jalr_id;
	wire lui_id;
	wire lbu_id;
	wire lhu_id;
	wire mfhi_id;
	wire mflo_id;
	wire mthi_id;
	wire mtlo_id;
	wire sb_id;
	wire sh_id;
	wire sign_sel_id;      // selector for sign or zero extend
	wire memWrite_id;//1-->active
	wire memRead_id; //1-active
	wire memToReg_id; // 0--> alu result   1--> memory data
	wire r31_select_id ;
	wire readenable_id; 
	wire [4:0] operation_id ;

      

	Control_unit  Control_unit (
		.opcode(opcode_id),
		.func(func_id),
		.sign_sel(sign_sel_id),
		.regDst(regDst_id),
		.aluSrc(aluSrc_id),
		.memRead(memRead_id),
		.memWrite(memWrite_id),
		.memToReg(memToReg_id),
		.readenable(readenable_id),
		.writeenable(regWrite_id),
		.beq(beq_id),
		.bne(bne_id),
		.blez(blez_id),
		.bgez(bgez_id),	
		.bgtz(bgtz_id),
		.jal(jal_id),
		.jr(jr_id),
		.j(j_id),
		.jalr(jalr_id),
		.r31_select(r31_select_id),
		.operation(operation_id),
		.lui(lui_id),
		.lbu(lbu_id),
		.lhu(lhu_id),
		.sh(sh_id),
		.sb(sb_id),
		.mfhi(mfhi_id),
		.mflo(mflo_id),	
		.mthi(mthi_id),
		.mtlo(mtlo_id)		
	);	
			


	//immediate extension 

	
	wire[31:0] sign_extended_id;
	reg[31:0] sign_extended16_id;
	
	integer i;
	
	always @(*)
		begin
		sign_extended16_id[15:0] <= instr_id[15:0];
		for (i=16; i<32;i=i+1)
		begin
			sign_extended16_id[i]<=instr_id[15];
		end
		end
		

	reg[31:0] zero_extended_id;
	
	always @(*)
		begin
		zero_extended_id[15:0] <= instr_id[15:0];
		for (i=12; i<32;i=i+1)
		begin
			zero_extended_id[i]<= 1'b0 ;
		end
		end
	
                                         	
	assign sign_extended_id =( sign_sel_id==1 )? sign_extended16_id : zero_extended_id;
	
	


	//====================================================== EX stage ================================================
	
	reg id_ex_reset;
	
	//instruction components
	reg[4:0]  rs_ex,rt_ex,rd_ex,shamt_ex;
	reg[31:0] sign_extended_ex;
	reg[25:0] jumpConst_ex;
	reg[5:0]  opcode_ex;
	reg[5:0]  func_ex;
	reg[31:0] pc_add_4_ex;
	reg[31:0] pc_add_1_ex;
	reg[15:0] imm16_ex;
	reg[31:0] lo_dataOut_ex;
	reg[31:0] hi_dataOut_ex;

	reg regWrite_ex;	//generated by control but not used now
	reg regDst_ex; 		//selector for the write register source (0--> rt or 1--> rd) 
	reg aluSrc_ex; 		//alu second operand source register 0--> from register file 1-->sign extended word
	reg memWrite_ex;	//1-->active
	reg memRead_ex; 	//1-active
	reg memToReg_ex; 	// 0--> alu result   1--> memory data
	reg [4:0] operation_ex;	
	reg beq_ex;
	reg bne_ex;
	reg blez_ex;
	reg bgez_ex;
	reg bgtz_ex;
	reg jal_ex;
	reg jr_ex;
	reg j_ex;
	reg jalr_ex;
	reg lui_ex;
	reg lbu_ex;
	reg lhu_ex;	
	reg r31_select_ex ;
	reg readenable_ex; 
	reg sb_ex;
	reg sh_ex;
	reg mfhi_ex;
	reg mflo_ex;
	reg mthi_ex;
	reg mtlo_ex;

	always @(posedge clk)
		begin
			if(id_ex_reset==1 || reset_b==0)
			begin
				regWrite_ex<=0;
				readenable_ex<=0;
				memWrite_ex<=0;
				memRead_ex<=0;
				beq_ex<=0;
				bne_ex<=0;
				blez_ex<=0;
				bgez_ex<=0;
				bgtz_ex<=0;
				jal_ex<=0;
				jr_ex<=0;
				j_ex<=0;
				jalr_ex<=0;
				lui_ex<=0;
				lbu_ex<=0;
				lhu_ex<=0;
				sb_ex<=0;
				sh_ex<=0;
				mfhi_ex<=0;
				mflo_ex<=0;
				mthi_ex<=0;
				mtlo_ex<=0;
				regDst_ex<=0; 
				operation_ex<=0;

			end
			else if(id_ex_enable==1)
			begin
				rs_ex<=rs_id;
				rt_ex<=rt_id;
				rd_ex<=rd_id;
				lo_dataOut_ex<=lo_dataOut_id;
				hi_dataOut_ex<=hi_dataOut_id;
				shamt_ex<=shamt_id;
				sign_extended_ex<=sign_extended_id;			
				regWrite_ex<=regWrite_id;
				regDst_ex<=regDst_id;
				r31_select_ex <= r31_select_id;
				aluSrc_ex<=aluSrc_id;
				beq_ex<=beq_id;
				bne_ex<=bne_id;
				blez_ex<=blez_id;
				bgez_ex<=bgez_id;
				bgtz_ex<=bgtz_id;
				jal_ex<=jal_id;
				jr_ex<=jr_id;
				j_ex<=j_id;
				jalr_ex<=jalr_id;
				lui_ex<=lui_id;
				lbu_ex<=lbu_id;
				lhu_ex<=lhu_id;
				mfhi_ex<=mfhi_id;
				mflo_ex<=mflo_id;
				mthi_ex<=mthi_id;
				mtlo_ex<=mtlo_id;
				memWrite_ex<=memWrite_id;
				memRead_ex<=memRead_id;
				memToReg_ex<=memToReg_id;
				readenable_ex<=readenable_id;	
				pc_add_4_ex<=pc_add_4_id;
				pc_add_1_ex<=pc_add_1_id; 
				jumpConst_ex<=jumpConst_id;
				operation_ex<=operation_id;
				opcode_ex<=opcode_id;
				func_ex<=func_id;
				imm16_ex<=imm16_id;
				sh_ex <= sh_id;
				sb_ex <= sb_id;
			end
		end
		
	 wire[4:0] rd_actual_ex;
	 wire[4:0]  rd_actual_ex1;
	 wire[4:0] R31=31;
	 assign rd_actual_ex1 = regDst_ex==0 ? rt_ex : rd_ex;
	 assign rd_actual_ex = r31_select_ex==0 ? rd_actual_ex1 : R31 ;
	 	 
	 
	 wire[31:0] aluOp1,aluOp2;
	 assign aluOp1=reg_rd1_ex;
	 assign aluOp2=aluSrc_ex ==0 ? reg_rd2_ex : sign_extended_ex;
	 
	 wire[31:0] aluResult_ex;
	 wire[31:0] aluResult_hi_ex;
	 wire aluZero_ex;
	 wire aluSign_ex;
	 
	 
	 ALU ALU
	 (
		.a(aluOp1),
		.b(aluOp2),
		.out_reg(aluResult_ex),
		.hi_out(aluResult_hi_ex),
		.shamt(shamt_ex),
		.zero_flag(aluZero_ex),
		.negative_flag(aluSign_ex),
		.operation(operation_ex)
	 );
	 
	 wire[31:0] pc_branch_ex , pc_jump_ex , pc_jumpr_ex ;
	 assign pc_branch_ex = (sign_extended_ex<<2)+pc_add_4_ex;
	 assign pc_jump_ex = { pc_add_4_ex[31:28] , (jumpConst_ex<<2) };
	 assign pc_jumpr_ex = reg_rd1_ex;
	
	 

	//============================================== MEM stage ================================================

	reg ex_mem_enable;
	reg ex_mem_reset;
	
	//instruction components
	reg [4:0] rs_mem,rt_mem;
	
	reg [4:0] rd_actual_mem;
	reg [31:0] reg_rd1_mem;	
	reg [31:0] reg_rd2_mem;
	reg [31:0] lo_dataOut_mem;
	reg [31:0] hi_dataOut_mem;

	reg[31:0] pc_add_4_mem;	

	reg aluZero_mem;
	reg aluSign_mem;
	reg[15:0] imm16_mem;
        reg[31:0] aluResult_mem;
	reg[31:0] aluResult_hi_mem; 
	
	reg regWrite_mem;
	reg beq_mem;
	reg bne_mem;
	reg blez_mem;
	reg bgez_mem;
	reg bgtz_mem;
	reg j_mem;
	reg jal_mem;
	reg jr_mem;
	reg jalr_mem;
	reg lui_mem;
	reg lbu_mem;
	reg lhu_mem;
	reg memWrite_mem;
	reg memRead_mem; 
	reg memToReg_mem;
	reg sb_mem;
	reg sh_mem;
	reg mfhi_mem;
	reg mflo_mem;
	reg mthi_mem;
	reg mtlo_mem;
	
	always @(posedge clk)
		begin
			if(ex_mem_reset==1 || reset_b==0)
			begin
				regWrite_mem<=0;
				beq_mem<=0;
				bne_mem<=0;
				blez_mem<=0;
				bgez_mem<=0;
				bgtz_mem<=0;
				j_mem<=0;
				jal_mem<=0;
				jr_mem<=0;
				jalr_mem<=0;
				memWrite_mem<=0;
				memRead_mem<=0;
				lui_mem<=0;
				lbu_mem<=0;
				lhu_mem<=0;
				sb_mem<=0;
				sh_mem<=0;
				mfhi_mem<=0;
				mflo_mem<=0;
				mthi_mem<=0;
				mtlo_mem<=0;
				memToReg_mem<=0;
			end
			if(ex_mem_enable==1)
			begin
				rs_mem<=rs_ex;
				rt_mem<=rt_ex;
				lo_dataOut_mem<=lo_dataOut_ex;
				hi_dataOut_mem<=hi_dataOut_ex;
				rd_actual_mem<=rd_actual_ex;
				reg_rd2_mem<=reg_rd2_ex;
				reg_rd1_mem<=reg_rd1_ex;
				aluResult_mem<=aluResult_ex;
				aluResult_hi_mem<=aluResult_hi_ex;
				aluZero_mem<=aluZero_ex;
				aluSign_mem<=aluSign_ex;
				beq_mem<=beq_ex;
				bne_mem<=bne_ex;
				blez_mem<=blez_ex;
				bgez_mem<=bgez_ex;
				bgtz_mem<=bgtz_ex;
				j_mem<=j_ex;
				jal_mem<=jal_ex;
				jr_mem<=jr_ex;
				jalr_mem<=jalr_ex;
				lui_mem<=lui_ex;
				lbu_mem<=lbu_ex;
				lhu_mem<=lhu_ex;
				mfhi_mem<=mfhi_ex;
				mflo_mem<=mflo_ex;
				mthi_mem<=mthi_ex;
				mtlo_mem<=mtlo_ex;
				pc_branch_mem<=pc_branch_ex;
				pc_jump_mem<=pc_jump_ex;
				pc_jumpr_mem<=pc_jumpr_ex;
				pc_add_4_mem<=pc_add_4_ex;
				sb_mem<=sb_ex;
				sh_mem<=sh_ex;
				regWrite_mem<=regWrite_ex;
				
				memWrite_mem<=memWrite_ex;
				memRead_mem<=memRead_ex;
				memToReg_mem<=memToReg_ex;
				imm16_mem<=imm16_ex;
			end
		end


	 assign beq_sel_mem=aluZero_mem & beq_mem;		
	 assign bne_sel_mem=( !aluZero_mem) & bne_mem; 
	 assign bgtz_sel_mem=( !aluSign_mem) & ( bgtz_mem);
	 assign blez_sel_mem=( aluZero_mem || aluSign_mem) & blez_mem;
	 assign bgez_sel_mem=( aluZero_mem || !aluSign_mem) & bgez_mem; 
	 assign jump_sel_mem=( j_mem || jal_mem );
	 assign jumpr_sel_mem=(jr_mem || jalr_mem );  
	 
	 
	 wire[31:0] mem_read_data_mem;
	 wire [31:0]  mem_wr_data_mem;	
 
	 DMem DM
	 (
		.address(aluResult_mem),
		.din(mem_wr_data_mem),
		.dout(mem_read_data_mem),
		.clk(clk),
		.read(memRead_mem),
		.write(memWrite_mem)
	 );

	wire[31:0] data_sh_in , data_sb_in;           // data written in memeory in sh and sb instr.
	assign data_sh_in = { reg_rd2_mem[15:0] , 16'b0 };
	assign data_sb_in = { reg_rd2_mem[7:0]  , 24'b0 };
	
	wire mem_wr_data_mem1;

	assign  mem_wr_data_mem1 = (sh_mem==1)? data_sh_in : reg_rd2_mem;
	assign  mem_wr_data_mem = (sb_mem==1)? data_sb_in : mem_wr_data_mem1;



	 //============================================== WB stage =================================================
	 
	 //instruction components
	reg[4:0] rs_wb,rt_wb;

	reg[31:0] pc_add_4_wb;	
        reg[31:0] reg_rd1_wb;
	reg jal_wb;	
	reg jalr_wb;
	reg lui_wb;
	reg lbu_wb;
	reg lhu_wb;
	reg mfhi_wb;
	reg mflo_wb;
	reg mthi_wb;
	reg mtlo_wb;
	reg[31:0] mem_read_data_wb;
	reg[31:0] aluResult_wb;
	reg[31:0] aluResult_hi_wb;
	reg[15:0] imm16_wb;

	reg[31:0] lo_dataOut_wb;
	reg[31:0] hi_dataOut_wb;

        reg memToReg_wb;
        wire[31:0] reg_wr_wb1;      // data in reg 
        wire[31:0] reg_wr_wb2;
        wire[31:0] reg_wr_wb3;
        wire[31:0] reg_wr_wb4;
        wire[31:0] reg_wr_wb5;
	wire[31:0] reg_wr_wb6;

	always @(posedge clk)
		begin
			if(reset_b==0)
			begin
				regWrite_wb<=0;
				memToReg_wb<=0;
				jal_wb<=0;
				jalr_wb<=0;
				lui_wb<=0;
				lbu_wb<=0;
				lhu_wb<=0;
				mfhi_wb<=0;
				mflo_wb<=0;
				mthi_wb<=0;
				mtlo_wb<=0;
			end
			else
			begin
				rs_wb<=rs_mem;
				rt_wb<=rt_mem;
				rd_actual_wb<=rd_actual_mem;
				reg_rd1_wb<= reg_rd1_mem;
				aluResult_wb<=aluResult_mem;
				aluResult_hi_wb<=aluResult_hi_mem;
				mem_read_data_wb<=mem_read_data_mem;
				imm16_wb<=imm16_mem;
				regWrite_wb<=regWrite_mem;
				memToReg_wb<=memToReg_mem;
				jal_wb<=jal_mem;
				jalr_wb<=jalr_mem;
				lui_wb<=lui_mem;
				lbu_wb<=lbu_mem;
				lhu_wb<=lhu_mem;
				mfhi_wb<=mfhi_mem;
				mflo_wb<=mflo_mem;
				mthi_wb<=mthi_mem;
				mtlo_wb<=mtlo_mem;				
				lo_dataOut_wb<=lo_dataOut_mem;
				hi_dataOut_wb<=hi_dataOut_mem;
				pc_add_4_wb<=pc_add_4_mem;
			end
			
		end

			wire[31:0] data_lui_wb;  // data written in lui instruction
			assign data_lui_wb = imm16_wb << 16 ;	
			
			wire[31:0] data_lhu_wb;
			assign data_lhu_wb = { 16'b0 , mem_read_data_wb[15:0] } ;
			
			wire[31:0] data_lbu_wb;
			assign data_lbu_wb = { 24'b0 , mem_read_data_wb[7:0] } ;	

		assign reg_wr_wb1 =memToReg_wb ==0 ? aluResult_wb : mem_read_data_wb;
		assign reg_wr_wb2 =( (jal_wb || jalr_wb )==0 )? reg_wr_wb1 : pc_add_4_wb;
		assign reg_wr_wb3 =(lui_wb==1)? data_lui_wb : reg_wr_wb2;
		assign reg_wr_wb4 =(lhu_wb==1)?  data_lhu_wb  : reg_wr_wb3;
		assign reg_wr_wb5 =(lbu_wb==1)?  data_lbu_wb  : reg_wr_wb4;
		assign reg_wr_wb6 =(mfhi_wb==1)?    hi_dataOut_wb   : reg_wr_wb5;
		assign reg_wr_wb  =(mflo_wb==1)?    lo_dataOut_wb   : reg_wr_wb6;

		 assign hi_dataIn_wb = (mthi_wb==1)? reg_rd1_wb : aluResult_hi_wb;
		 assign lo_dataIn_wb = (mtlo_wb==1)? reg_rd1_wb : aluResult_wb; 

	//======================================= Hazard ===============================================
	
	
	//stall control outputs:
	//pc_en_id
	//if_id_enable
	//id_ex_enable
	//ex_mem_enable
	
	wire data_hazard;
	
	assign data_hazard= /*ex-id hazards*/ ( (rs_id==rd_actual_ex) && (regWrite_ex==1) ) ||
			((rt_id==rd_actual_ex) && (regWrite_ex==1) ) ||
			/*mem-id hazards*/ ( (rs_id==rd_actual_mem) && (regWrite_mem==1) )||
			( (rt_id==rd_actual_mem) && (regWrite_mem==1) );
			
	wire control_hazard;
	assign control_hazard= (beq_mem==1 && aluZero_mem==1) || 
			( bne_mem==1 && aluZero_mem==0 ) ||
			( (bgtz_mem==1) && aluSign_mem==0 ) ||
			( blez_mem==1 && (aluZero_mem==1 || aluSign_mem==1) ) ||
			( bgez_mem==1 && (aluZero_mem==1 || aluSign_mem==0) ) || 
			( j_mem==1) || (jal_mem==1) || (jr_mem==1) || (jalr_mem==1) ;   
	
	always @(*)
	begin
		pc_en_id=1;
		lo_en_id= (mflo_id==1 || mtlo_id==1 || func_id==6'b011010 || func_id==6'b011011 || func_id==6'b011000 || func_id==6'b011001)? 1 : 0 ;
		hi_en_id= (mfhi_id==1 || mthi_id==1 || func_id==6'b011010 || func_id==6'b011011 || func_id==6'b011000 || func_id==6'b011001)? 1 : 0 ;
		if_id_enable=1;
		id_ex_enable=1;
		
		ex_mem_enable=1;
		
		id_ex_reset=0;
		ex_mem_reset=0;
		

		
		//r-instruction hazards
		if(data_hazard)
			begin
				pc_en_id=0;
				if_id_enable=0;
				id_ex_reset=1;
			end
		//control hazards (predict not taken)
		if(control_hazard)
		begin
			pc_en_id=1;
			id_ex_reset=1;
			ex_mem_reset=1;
		end
	end
endmodule
